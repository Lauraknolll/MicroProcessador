library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM_instrucoes is
   port( 
        clk      : in std_logic;
        endereco : in unsigned(6 downto 0);
        dado     : out unsigned(15 downto 0) 
   );
end entity;

architecture a_ROM_instrucoes of ROM_instrucoes is
   type mem is array (0 to 127) of unsigned(15 downto 0);
   constant conteudo_rom : mem := (
      -- caso endereco => conteudo
      --MOV destino, fonte

      0   => "0010000000010100", --ADDI A, 20
      1   => "0011000000000101", --SUBI A, 5
      2   => "1100000000000010", --LD R0, 2
      3   => "0100000000000000", --ADD A, R0
      4   => "1101100000001010", --LD B, 10
      5   => "0101100010000000", --SUB B, R1        
      6   => "0110100010000000", --AND B, R1
      7   => "0111000000000000", --OR A, R0
      8   => "1101100000001000", --LD B, 8
      9   => "1100001101000000", --LD R3, 64
      10  => "1110100100000000", --MOV B, R2
      11  => "1110000001000000", --MOV R0, A
      12  => "1101000000100000", --LD A, 32 
      13  => "1001000110000000", --COMP A,R3
      14  => "1011100000001111", --BHI  +15    -- EH PARA FALHAR A < R3
      15  => "1001000100000000", --COMP A, R2
      16  => "1011100000000011", --BHI +3       --VAI DAR CERTO

      17  => "1001011100110011", --NOP         --EH PARA FALHAR
      18  => "1111000000110010", --JUMP 50     --EH PARA FALHAR
      
      19  => "1001100000000000",  --COMP B, R0
      20  => "1010000111110110",  -- BGE -10   --EH PARA FALHAR
      21  => "1100010000001000",  -- LD R4,8
      22  => "1001101000000000",  -- COMP B, R4
      23  => "1010000000000101",  -- BGE +5   -- VAI DAR CERTO

      24  => "1111110001000000",  -- JUMP 64
      25  => "1001011100110011",  --NOP
      26  => "1001011100110011",  --NOP
      27  => "1001011100110011",  --NOP
      28  => "1001011100110011",  --NOP

      29  => "1100101000001000",  --LD R10, 8
      30  => "1101100000100000",  --LD B, 32
      31  => "1000000000000000",  --SW
      32  => "1101100000000000",  --LD B, 0
      33  => "0001000000000000",  -- LW -- O VALOR ESTARÁ NO ACC B
      34  => "0000000000000000",  -- EXCEÇÃO
      -- 35  => "1110010101000000",  --
      -- 36  => "1110001100000000",  --
      -- 37  => "0100001100000000",  --
      -- 38  => "1001001000000000",  --
      -- 39  => "1010000000000100",  -- 
      -- 40  => "1110010100000000",  --
      -- 41  => "1000000000000000",  --
      -- 42  => "1111000000100101",  --JUMP 
      -- 43  => "1110001011000000",  --MOV A, R5
      -- 44  => "1110010100000000",  --MOV R10, A
      -- 45  => "1111000000010110",  --JUMP 
      -- 46  => "1001011100110011",  --NOP

      -- --Leitura dos números primos até 1024
      -- 47  => "1100101000000010",  --LD R10, 2
      -- 48  => "1101000000000000",  --LD A, 0
      -- 49  => "1101100000000001",  --LD B, 0
      -- 50  => "1110010101000000",  --MOV A, R10

      -- 51  => "1001001000000000",  --COMP A, R4 
      -- 52  => "1010000000001011",  --BGE 
      -- 53  => "0001000000000000",  --LW
      -- 54  => "1001100100000000",  --COMP B, R2
      -- 55  => "1010000000000010",  --BGE
      -- 56  => "1111000000111011",  --JUMP 
      -- 57  => "1110010101000000",  --MOV A, R10
      -- 58  => "1110000000000000",  --MOV R0, A
      -- 59  => "1110010101000000",  --MOV A, R10   
      -- 60  => "0010000000000001",  --ADDI A, 1
      -- 61  => "1110010100000000",  --MOV R10, A
      -- 62  => "1111000000110011",  --JUMP  

      -- 63  => "1001011100110011",  --NOP
      -- 64  => "0000000000000000", --EXCEÇÃO
      -- 65  => "1001011100110011",  --NOP
      -- abaixo: casos omissos => (zero em todos os bits)
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;