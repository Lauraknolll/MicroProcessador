library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TopLevel is
    port (
        clock : in std_logic;
        dado_escrita_banco : in unsigned(15 downto 0);
        reset_b, reset_acc : in std_logic; --o reset dos dois acumuladores é o mesmo??
        qual_reg_escreve, qual_reg_le : in unsigned(3 downto 0); --no banco
        escreve_banco : in std_logic;

        escolhe_accA, escolhe_accB : in std_logic; 
        dado_escrita_acc : in unsigned(15 downto 0);

        op_com_cte : in std_logic; --se for 1 é ADDI ou SUBI 
        cte : in unsigned(15 downto 0); --a cte que vem da instrução

        sel0, sel1 : in std_logic; --operações da ula
        carry, overflow, zero, sinal : out std_logic;
        --descobrir quais as entradas e saídas que precisa

        op_mov_p_reg, op_mov_p_acc, op_ld_acc : in std_logic
    );
end entity;

architecture struct of TopLevel is

    component reg16bits is
        port( 
            clk      : in std_logic;
            rst      : in std_logic;
            wr_en    : in std_logic;
            data_in  : in unsigned(15 downto 0);
            data_out : out unsigned(15 downto 0)
        );
    end component;

    component BancoReg is
        port( 
            clk_b         : in std_logic;
            rst_b          : in std_logic; 
            wr_en         : in std_logic; 
            sel_reg_wr    : in unsigned(3 downto 0); 
            sel_reg_rd    : in unsigned(3 downto 0); 
            --acc           : in std_logic; 
            data_wr       : in unsigned(15 downto 0); 
            data_out_r1   : out unsigned(15 downto 0) 
        );
    end component;

    component ULA is
        port(
            in_A, in_B : in unsigned(15 downto 0);
            Sel0, Sel1 : in std_logic;
            Resultado : out unsigned(15 downto 0);
            Carry, Overflow, Zero, Sinal : out std_logic
        );
    end component;

    signal banco_ula, ula_accs, acc0_ula, acc1_ula, accs_ula, dado_ula, escrita_banco, escrita_acc : unsigned(15 downto 0);
    signal escolhe_acc1 : std_logic;

begin

    --MUX entrada do banco
    escrita_banco <= dado_escrita_banco when op_mov_p_reg = '0' else --quando é LD em algum reg
                    accs_ula when op_mov_p_reg = '1' else --quando é MOV acc, reg
                    (others => '0');

    uut0 : BancoReg port map (clk_b => clock, rst_b => reset_b, wr_en => escreve_banco, sel_reg_wr => qual_reg_escreve, sel_reg_rd => qual_reg_le, data_wr => escrita_banco, data_out_r1 => banco_ula);
    --MUX entrada dos acumuladores A e B
    escrita_acc <= banco_ula when (op_mov_p_acc = '1' and op_ld_acc = '0') else
                    dado_escrita_acc when (op_mov_p_acc = '0' and op_ld_acc = '1') else
                    ula_accs when (op_mov_p_acc = '0' and op_ld_acc = '0') else
                    (others => '0');
                    
    uutA : reg16bits port map (clk => clock, rst => reset_acc, wr_en => escolhe_accA, data_in => escrita_acc, data_out => acc0_ula); --acumulador A/0

    uutB : reg16bits port map (clk => clock, rst => reset_acc, wr_en => escolhe_accB, data_in => escrita_acc, data_out => acc1_ula); --acumulador B/1
    --MUX da saída do banco e da cte na entrada A da ula
    dado_ula <= banco_ula when op_com_cte = '0' else
                cte when op_com_cte = '1' else
                (others => '0');
    --MUX da saída dos acc na entrada B da ula
    accs_ula <= acc0_ula when escolhe_accA = '1' else
                acc1_ula when escolhe_accB = '1' else
                (others => '0');
    uut1 : ULA port map (in_A => dado_ula, in_B => accs_ula, Sel0 => sel0, Sel1 => sel1, Resultado => ula_accs, Carry => carry, Overflow => overflow, Zero => zero, Sinal => sinal);

end struct ; 