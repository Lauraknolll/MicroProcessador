library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
   port( 
        clk      : in std_logic;
        endereco : in unsigned(6 downto 0);
        dado     : out unsigned(15 downto 0) 
   );
end entity;

architecture a_ROM of ROM is
   type mem is array (0 to 127) of unsigned(15 downto 0);
   constant conteudo_rom : mem := (
      -- caso endereco => conteudo
      --MOV destino, fonte

      --Colocar o 1024 no R4
      0   => "1101000001111111", --LD A, 127
      1   => "0010000000000001", --ADDI A, 1
      2   => "1110001000000000", --MOV R4, A
      3   => "0100001000000000", --ADD A, R4
      4   => "1110001000000000", --MOV R4, A
      5   => "0100001000000000", --ADD A, R4        
      6   => "1110001000000000", --MOV R4, A
      7   => "0100001000000000", --ADD A, R4
      8   => "1110001000000000", --MOV R4, A
      
      --Colocar 1 em todas as posições de 0 a 1023
      9   => "1100101000000000", --LD R10, 0
      10  => "1101100000000001", --LD B, 1
      11  => "1110010101000000", --MOV A, R10
      12  => "1001001000000000", --COMP A, R4 
      13  => "1010000000000110", --BGE 
      14  => "1000000000000000", --SW 
      15  => "0100110100000000", --ADD B, R10
      16  => "1110110100000000", --MOV R10, B
      17  => "1101100000000001", --LD B, 1
      18  => "1111000000001011", --JUMP

      --Crivo de Erastóteles
      19  => "1100001000000001",  --LD R2, 1
      20  => "1100101000000010",  --LD R10, 2
      21  => "1100001100100001",  --LD R3, 33
      22  => "1110010101000000",  --MOV A, R10
      23  => "1001000110000000",  --COMP A, R3
      24  => "1010000000010110",  --BGE 
      25  => "0001000000000000",  --LW
      26  => "1110110010000000",  --MOV R9, B
      27  => "1110110101000000",  --MOV B, R10
      28  => "0010100000000001",  --ADDI B, 1
      29  => "1110101010000000",  --MOV R5, B
      30  => "1110010011000000",  --MOV A, R9
      31  => "1001000100000000",  --COMP A, R2
      32  => "1010000000000010",  --BGE 
      33  => "1111000000101011",  --JUMP 
      34  => "1101100000000000",  --LD B, 0
      35  => "1110010101000000",  --MOV A, R10
      36  => "1110001100000000",  --MOV R6, A
      37  => "0100001100000000",  --ADD A, R6
      38  => "1001001000000000",  --COMP A, R4
      39  => "1010000000000100",  --BGE 
      40  => "1110010100000000",  --MOV R10, A
      41  => "1000000000000000",  --SW
      42  => "1111000000100101",  --JUMP 
      43  => "1110001011000000",  --MOV A, R5
      44  => "1110010100000000",  --MOV R10, A
      45  => "1111000000010110",  --JUMP 
      46  => "1001011100110011",  --NOP

      --Leitura dos números primos até 1024
      47  => "1100101000000010",  --LD R10, 2
      48  => "1101000000000000",  --LD A, 0
      49  => "1101100000000001",  --LD B, 0
      50  => "1110010101000000",  --MOV A, R10

      51  => "1001001000000000",  --COMP A, R4 
      52  => "1010000000001011",  --BGE 
      53  => "0001000000000000",  --LW
      54  => "1001100100000000",  --COMP B, R2
      55  => "1010000000000010",  --BGE
      56  => "1111000000111011",  --JUMP 
      57  => "1110010101000000",  --MOV A, R10
      58  => "1110000000000000",  --MOV R0, A
      59  => "1110010101000000",  --MOV A, R10   
      60  => "0010000000000001",  --ADDI A, 1
      61  => "1110010100000000",  --MOV R10, A
      62  => "1111000000110011",  --JUMP  

      63  => "1001011100110011",  --NOP
      64  => "0000000000000000", --EXCEÇÃO
      65  => "1001011100110011",  --NOP
      -- abaixo: casos omissos => (zero em todos os bits)
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;