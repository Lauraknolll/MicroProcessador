library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
   port( 
        clk      : in std_logic;
        endereco : in unsigned(6 downto 0);
        dado     : out unsigned(15 downto 0) 
   );
end entity;

architecture a_ROM of ROM is
   type mem is array (0 to 127) of unsigned(15 downto 0);
   constant conteudo_rom : mem := (
      -- caso endereco => conteudo
      --MOV destino, fonte

      -- TESTE DE TODAS AS INSTRUÇÕES -------------------------

      0   => "0010000000010100", --ADDI A, 20
      1   => "0011000000000101", --SUBI A, 5
      2   => "1100000000000010", --LD R0, 2
      3   => "0100000000000000", --ADD A, R0
      4   => "1101100000001010", --LD B, 10
      5   => "0101100000000000", --SUB B, R0        
      6   => "0110100000000000", --AND B, R0         
      7   => "0111000000000000", --OR A, R0        
      8   => "1101100000001000", --LD B, 8
      9   => "1100001101000000", --LD R3, 64
      10  => "1100001000000111", --LD R2, 7
      11  => "1110100101000000", --MOV B, R2   
      12  => "1110000001000000", --MOV R0, A   
      13  => "1101000000100000", --LD A, 32 
      14  => "1001000110000000", --COMP A,R3
      15  => "1011100000001111", --BHI  
      16  => "1001000100000000", --COMP A, R2
      17  => "1011100000000011", --BHI 

      18  => "1001011100110011", --NOP         
      19  => "1111000000110010", --JUMP 50     
      
      20  => "1001100110000000", --COMP B, R3
      21  => "1010000111110110", --BGE -10  
      22  => "1100010000000111", --LD R4,7
      23  => "1001101000000000", --COMP B, R4
      24  => "1010000000000101", --BGE  

      25  => "1111110001000000", --JUMP 64
      26  => "1001011100110011", --NOP
      27  => "1001011100110011", --NOP
      28  => "1001011100110011", --NOP
      
      29  => "1001011100110011", --NOP
      30  => "1100101000001000", --LD R10, 8
      31  => "1101100000100000", --LD B, 32
      32  => "1111000001000000", --JUMP 64

      64  => "1000000000000000", --SW
      65  => "1101100000000000", --LD B, 0
      66  => "0001000000000000", --LW 
      67  => "0000000000000000", --EXCEÇÃO


      -- VALIDAÇÃOOOOOOOO -------------------------------

      --Colocar o 1024 no R4
      -- 0   => "1101000001111111", --LD A, 127
      -- 1   => "0010000000000001", --ADDI A, 1
      -- 2   => "1110001000000000", --MOV R4, A
      -- 3   => "0100001000000000", --ADD A, R4
      -- 4   => "1110001000000000", --MOV R4, A
      -- 5   => "0100001000000000", --ADD A, R4        
      -- 6   => "1110001000000000", --MOV R4, A
      -- 7   => "0100001000000000", --ADD A, R4
      -- 8   => "1110001000000000", --MOV R4, A
      
      -- --Colocar 1 em todas as posições de 0 a 1023
      -- 9   => "1100101000000000", --LD R10, 0
      -- 10  => "1101100000000001", --LD B, 1
      -- 11  => "1110010101000000", --MOV A, R10
      -- 12  => "1001001000000000", --COMP A, R4 
      -- 13  => "1010000000000110", --BGE 
      -- 14  => "1000000000000000", --SW 
      -- 15  => "0100110100000000", --ADD B, R10
      -- 16  => "1110110100000000", --MOV R10, B
      -- 17  => "1101100000000001", --LD B, 1
      -- 18  => "1111000000001011", --JUMP

      -- --Crivo de Erastóteles
      -- 19  => "1100001000000001",  --LD R2, 1
      -- 20  => "1100101000000010",  --LD R10, 2
      -- 21  => "1100001100100001",  --LD R3, 33
      -- 22  => "1110010101000000",  --MOV A, R10
      -- 23  => "1001000110000000",  --COMP A, R3
      -- 24  => "1010000000010110",  --BGE 
      -- 25  => "0001000000000000",  --LW
      -- 26  => "1110110010000000",  --MOV R9, B
      -- 27  => "1110110101000000",  --MOV B, R10
      -- 28  => "0010100000000001",  --ADDI B, 1
      -- 29  => "1110101010000000",  --MOV R5, B
      -- 30  => "1110010011000000",  --MOV A, R9
      -- 31  => "1001000100000000",  --COMP A, R2
      -- 32  => "1010000000000010",  --BGE 
      -- 33  => "1111000000101011",  --JUMP 
      -- 34  => "1101100000000000",  --LD B, 0
      -- 35  => "1110010101000000",  --MOV A, R10
      -- 36  => "1110001100000000",  --MOV R6, A
      -- 37  => "0100001100000000",  --ADD A, R6
      -- 38  => "1001001000000000",  --COMP A, R4
      -- 39  => "1010000000000100",  --BGE 
      -- 40  => "1110010100000000",  --MOV R10, A
      -- 41  => "1000000000000000",  --SW
      -- 42  => "1111000000100101",  --JUMP 
      -- 43  => "1110001011000000",  --MOV A, R5
      -- 44  => "1110010100000000",  --MOV R10, A
      -- 45  => "1111000000010110",  --JUMP 
      -- 46  => "1001011100110011",  --NOP

      -- --Leitura dos números primos até 1024
      -- 47  => "1100101000000010",  --LD R10, 2
      -- 48  => "1101000000000000",  --LD A, 0
      -- 49  => "1101100000000001",  --LD B, 0
      -- 50  => "1110010101000000",  --MOV A, R10

      -- 51  => "1001001000000000",  --COMP A, R4 
      -- 52  => "1010000000001011",  --BGE 
      -- 53  => "0001000000000000",  --LW
      -- 54  => "1001100100000000",  --COMP B, R2
      -- 55  => "1010000000000010",  --BGE
      -- 56  => "1111000000111011",  --JUMP 
      -- 57  => "1110010101000000",  --MOV A, R10
      -- 58  => "1110000000000000",  --MOV R0, A
      -- 59  => "1110010101000000",  --MOV A, R10   
      -- 60  => "0010000000000001",  --ADDI A, 1
      -- 61  => "1110010100000000",  --MOV R10, A
      -- 62  => "1111000000110011",  --JUMP  

      -- 63  => "1001011100110011",  --NOP
      -- 64  => "0000000000000000", --EXCEÇÃO
      -- 65  => "1001011100110011",  --NOP

      -- -- abaixo: casos omissos => (zero em todos os bits)
      others => (others=>'0')
   );
begin
   process(clk)
   begin
      if(rising_edge(clk)) then
         dado <= conteudo_rom(to_integer(endereco));
      end if;
   end process;
end architecture;